module mul32 #(parameter T = 0.000, parameter N = 32)(
    input [N-1:0] a,
    input [N-1:0] b,
    input mode,
    output [N-1:0] hi,
    output [N-1:0] lo
);
    // Error is in bits: 48, 47, 46, 45
    wire c;
    wire c_;
    wire prod_comp;
    wire [N-1:0] a_;
    wire [N-1:0] b_;
    wire [N-1:0] a__;
    wire [N-1:0] b__;
    wire [N-1:0] lo_;
    wire [N-1:0] hi_;
    wire [N-1:0] lo__;
    wire [N-1:0] hi__;
    wire [N-1:0] s0 [2*N-2:0];
    wire [N-1:0] s1 [2*N-2:0];
    wire [N-1:0] s2 [2*N-2:0];
    wire [N-1:0] s3 [2*N-2:0];
    wire [N-1:0] s4 [2*N-2:0];
    wire [N-1:0] s5 [2*N-2:0];
    wire [N-1:0] s6 [2*N-2:0];
    wire [N-1:0] s7 [2*N-2:0];
    wire [N-1:0] s8 [2*N-2:0];
    genvar w;
    genvar j;
    genvar k;

    assign a_ = a^{(N-1){mode&a[N-1]}};
    assign b_ = b^{(N-1){mode&b[N-1]}};
    assign prod_comp = a[N-1]^b[N-1];
    assign lo__ = lo_^{(N-1){prod_comp}};
    assign hi__ = hi_^{(N-1){prod_comp}};
    add32 #(.T(T)) a_comp(
        .a(a_),
        .b(32'h00000000),
        .c_1(a[N-1]),
        .s(a__)
    );
    add32 #(.T(T)) b_comp(
        .a(b_),
        .b(32'h00000000),
        .c_1(b[N-1]),
        .s(b__)
    );

    generate
        // Stage 0: Partial-products generation
        for(w = 0;w <= 2*N-2;w = w+1)
        begin
            if(w < N)
            begin
                for(j = 0;j <= w;j = j+1)
                    assign #(T) s0[w][j] = a__[w-j]&b__[j];
                // for(k = w+1;k < N;k = k+1)
                //     assign s0[w][k] = 1'b0;
            end
            else
            begin
                for(j = 0;j < 2*N - 1 - w;j = j+1)
                    assign #(T) s0[w][j] = a__[N-1-j]&b__[w+j+1-N];
                // for(k = 2*N-w;k < N;k = k+1)
                //     assign s0[w][k] = 1'b0;
            end
        end
        // Stage 1
        // Max depth: 28 (27:0)
        for(w = 0;w <= 2*N-2;w = w+1)
        begin
            case(w)
                28:
                begin
                    ha #(.T(T)) ha1(.i(s0[w][1:0]),.o({s1[w+1][0],s1[w][0]}));
                    assign s1[w][27:1] = s0[w][28:2];
                end
                29:
                begin
                    fa #(.T(T)) fa1(.i(s0[w][2:0]),.o({s1[w+1][0],s1[w][1]}));
                    ha #(.T(T)) ha2(.i(s0[w][4:3]),.o({s1[w+1][1],s1[w][2]}));
                    assign s1[w][27:3] = s0[w][29:5];
                end
                30:
                begin
                    fa #(.T(T)) fa2(.i(s0[w][2:0]),.o({s1[w+1][0],s1[w][2]}));
                    fa #(.T(T)) fa3(.i(s0[w][5:3]),.o({s1[w+1][1],s1[w][3]}));
                    ha #(.T(T)) ha3(.i(s0[w][7:6]),.o({s1[w+1][2],s1[w][4]}));
                    assign s1[w][27:5] = s0[w][30:8];
                end
                31:
                begin
                    fa #(.T(T)) fa4(.i(s0[w][2:0]),.o({s1[w+1][0],s1[w][3]}));
                    fa #(.T(T)) fa5(.i(s0[w][5:3]),.o({s1[w+1][1],s1[w][4]}));
                    fa #(.T(T)) fa6(.i(s0[w][8:6]),.o({s1[w+1][2],s1[w][5]}));
                    ha #(.T(T)) ha4(.i(s0[w][10:9]),.o({s1[w+1][3],s1[w][6]}));
                    assign s1[w][27:7] = s0[w][31:11];
                end
                32:
                begin
                    fa #(.T(T)) fa7(.i(s0[w][2:0]),.o({s1[w+1][0],s1[w][4]}));
                    fa #(.T(T)) fa8(.i(s0[w][5:3]),.o({s1[w+1][1],s1[w][5]}));
                    fa #(.T(T)) fa9(.i(s0[w][8:6]),.o({s1[w+1][2],s1[w][6]}));
                    ha #(.T(T)) ha5(.i(s0[w][10:9]),.o({s1[w+1][3],s1[w][7]}));
                    assign s1[w][27:8] = s0[w][30:11];
                end
                33:
                begin
                    fa #(.T(T)) fa10(.i(s0[w][2:0]),.o({s1[w+1][0],s1[w][4]}));
                    fa #(.T(T)) fa11(.i(s0[w][5:3]),.o({s1[w+1][1],s1[w][5]}));
                    fa #(.T(T)) fa12(.i(s0[w][8:6]),.o({s1[w+1][2],s1[w][6]}));
                    assign s1[w][27:7] = s0[w][29:9];
                end
                34:
                begin
                    fa #(.T(T)) fa13(.i(s0[w][2:0]),.o({s1[w+1][0],s1[w][3]}));
                    fa #(.T(T)) fa14(.i(s0[w][5:3]),.o({s1[w+1][1],s1[w][4]}));
                    assign s1[w][27:5] = s0[w][28:6];
                end
                35:
                begin
                    fa #(.T(T)) fa15(.i(s0[w][2:0]),.o({s1[w+1][0],s1[w][2]}));
                    assign s1[w][27:3] = s0[w][27:3];
                end
                36:
                begin
                    assign s1[w][27:1] = s0[w][26:0];
                end
                default:
                    assign s1[w] = s0[w];
            endcase 
        end
        // Stage 2
        // Max depth: 19 (18:0)
        for(w = 0;w <= 2*N-2;w = w+1)
        begin
            case(w)
                19:
                begin
                    // fa - 0, ha - 1
                    ha #(.T(T)) ha1(.i(s1[w][1:0]),.o({s2[w+1][0],s2[w][0]}));
                    assign s2[w][18:1] = s1[w][19:2];
                end
                20:
                begin
                    // fa - 1, ha - 1
                    fa #(.T(T)) fa1(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][1]}));
                    ha #(.T(T)) ha2(.i(s1[w][4:3]),.o({s2[w+1][1],s2[w][2]}));
                    assign s2[w][18:3] = s1[w][20:5];
                end
                21:
                begin
                    // fa - 2, ha - 1
                    fa #(.T(T)) fa2(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][2]}));
                    fa #(.T(T)) fa3(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][3]}));
                    ha #(.T(T)) ha3(.i(s1[w][7:6]),.o({s2[w+1][2],s2[w][4]}));
                    assign s2[w][18:5] = s1[w][21:8];
                end
                22:
                begin
                    // fa - 3, ha - 1
                    fa #(.T(T)) fa4(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][3]}));
                    fa #(.T(T)) fa5(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][4]}));
                    fa #(.T(T)) fa6(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][5]}));
                    ha #(.T(T)) ha4(.i(s1[w][10:9]),.o({s2[w+1][3],s2[w][6]}));
                    assign s2[w][18:7] = s1[w][22:11];
                end
                23:
                begin
                    // fa - 4, ha - 1
                    fa #(.T(T)) fa7(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][4]}));
                    fa #(.T(T)) fa8(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][5]}));
                    fa #(.T(T)) fa9(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][6]}));
                    fa #(.T(T)) fa10(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][7]}));
                    ha #(.T(T)) ha5(.i(s1[w][13:12]),.o({s2[w+1][4],s2[w][8]}));
                    assign s2[w][18:9] = s1[w][23:14];
                end
                24:
                begin
                    // fa - 5, ha - 1
                    fa #(.T(T)) fa11(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][5]}));
                    fa #(.T(T)) fa12(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][6]}));
                    fa #(.T(T)) fa13(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][7]}));
                    fa #(.T(T)) fa14(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][8]}));
                    fa #(.T(T)) fa15(.i(s1[w][14:12]),.o({s2[w+1][4],s2[w][9]}));
                    ha #(.T(T)) ha6(.i(s1[w][16:15]),.o({s2[w+1][5],s2[w][10]}));
                    assign s2[w][18:11] = s1[w][24:17];
                end
                25:
                begin
                    // fa - 6, ha - 1
                    fa #(.T(T)) fa16(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][6]}));
                    fa #(.T(T)) fa17(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][7]}));
                    fa #(.T(T)) fa18(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][8]}));
                    fa #(.T(T)) fa19(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][9]}));
                    fa #(.T(T)) fa20(.i(s1[w][14:12]),.o({s2[w+1][4],s2[w][10]}));
                    fa #(.T(T)) fa21(.i(s1[w][17:15]),.o({s2[w+1][5],s2[w][11]}));
                    ha #(.T(T)) ha7(.i(s1[w][19:18]),.o({s2[w+1][6],s2[w][12]}));
                    assign s2[w][18:13] = s1[w][25:20];
                end
                26:
                begin
                    // fa - 7, ha - 1
                    fa #(.T(T)) fa22(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][7]}));
                    fa #(.T(T)) fa23(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][8]}));
                    fa #(.T(T)) fa24(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][9]}));
                    fa #(.T(T)) fa25(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][10]}));
                    fa #(.T(T)) fa26(.i(s1[w][14:12]),.o({s2[w+1][4],s2[w][11]}));
                    fa #(.T(T)) fa27(.i(s1[w][17:15]),.o({s2[w+1][5],s2[w][12]}));
                    fa #(.T(T)) fa28(.i(s1[w][20:18]),.o({s2[w+1][6],s2[w][13]}));
                    ha #(.T(T)) ha8(.i(s1[w][22:21]),.o({s2[w+1][7],s2[w][14]}));
                    assign s2[w][18:15] = s1[w][26:23];
                end
                27:
                begin
                    // fa - 8, ha - 1
                    fa #(.T(T)) fa29(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][8]}));
                    fa #(.T(T)) fa30(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][9]}));
                    fa #(.T(T)) fa31(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][10]}));
                    fa #(.T(T)) fa32(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][11]}));
                    fa #(.T(T)) fa33(.i(s1[w][14:12]),.o({s2[w+1][4],s2[w][12]}));
                    fa #(.T(T)) fa34(.i(s1[w][17:15]),.o({s2[w+1][5],s2[w][13]}));
                    fa #(.T(T)) fa35(.i(s1[w][20:18]),.o({s2[w+1][6],s2[w][14]}));
                    fa #(.T(T)) fa36(.i(s1[w][23:21]),.o({s2[w+1][7],s2[w][15]}));
                    ha #(.T(T)) ha9(.i(s1[w][25:24]),.o({s2[w+1][8],s2[w][16]}));
                    assign s2[w][18:17] = s1[w][27:26];
                end
                28, 29, 30, 31, 32, 33, 34, 35, 36:
                begin
                    // fa - 9, ha - 0
                    fa #(.T(T)) fa37(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][9]}));
                    fa #(.T(T)) fa38(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][10]}));
                    fa #(.T(T)) fa39(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][11]}));
                    fa #(.T(T)) fa40(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][12]}));
                    fa #(.T(T)) fa41(.i(s1[w][14:12]),.o({s2[w+1][4],s2[w][13]}));
                    fa #(.T(T)) fa42(.i(s1[w][17:15]),.o({s2[w+1][5],s2[w][14]}));
                    fa #(.T(T)) fa43(.i(s1[w][20:18]),.o({s2[w+1][6],s2[w][15]}));
                    fa #(.T(T)) fa44(.i(s1[w][23:21]),.o({s2[w+1][7],s2[w][16]}));
                    fa #(.T(T)) fa45(.i(s1[w][26:24]),.o({s2[w+1][8],s2[w][17]}));
                    assign s2[w][18] = s1[w][27];
                end
                37:
                begin
                    // fa - 8, ha - 0
                    fa #(.T(T)) fa46(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][9]}));
                    fa #(.T(T)) fa47(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][10]}));
                    fa #(.T(T)) fa48(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][11]}));
                    fa #(.T(T)) fa49(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][12]}));
                    fa #(.T(T)) fa50(.i(s1[w][14:12]),.o({s2[w+1][4],s2[w][13]}));
                    fa #(.T(T)) fa51(.i(s1[w][17:15]),.o({s2[w+1][5],s2[w][14]}));
                    fa #(.T(T)) fa52(.i(s1[w][20:18]),.o({s2[w+1][6],s2[w][15]}));
                    fa #(.T(T)) fa53(.i(s1[w][23:21]),.o({s2[w+1][7],s2[w][16]}));
                    assign s2[w][18:17] = s1[w][25:24];
                end
                38:
                begin
                    // fa - 7, ha - 0
                    fa #(.T(T)) fa54(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][8]}));
                    fa #(.T(T)) fa55(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][9]}));
                    fa #(.T(T)) fa56(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][10]}));
                    fa #(.T(T)) fa57(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][11]}));
                    fa #(.T(T)) fa58(.i(s1[w][14:12]),.o({s2[w+1][4],s2[w][12]}));
                    fa #(.T(T)) fa59(.i(s1[w][17:15]),.o({s2[w+1][5],s2[w][13]}));
                    fa #(.T(T)) fa60(.i(s1[w][20:18]),.o({s2[w+1][6],s2[w][14]}));
                    assign s2[w][18:15] = s1[w][24:21];
                end
                39:
                begin
                    // fa - 6, ha - 0
                    fa #(.T(T)) fa61(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][7]}));
                    fa #(.T(T)) fa62(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][8]}));
                    fa #(.T(T)) fa63(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][9]}));
                    fa #(.T(T)) fa64(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][10]}));
                    fa #(.T(T)) fa65(.i(s1[w][14:12]),.o({s2[w+1][4],s2[w][11]}));
                    fa #(.T(T)) fa66(.i(s1[w][17:15]),.o({s2[w+1][5],s2[w][12]}));
                    assign s2[w][18:13] = s1[w][23:18];
                end
                40:
                begin
                    // fa - 5, ha - 0
                    fa #(.T(T)) fa67(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][6]}));
                    fa #(.T(T)) fa68(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][7]}));
                    fa #(.T(T)) fa69(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][8]}));
                    fa #(.T(T)) fa70(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][9]}));
                    fa #(.T(T)) fa71(.i(s1[w][14:12]),.o({s2[w+1][4],s2[w][10]}));
                    assign s2[w][18:11] = s1[w][22:15];
                end
                41:
                begin
                    // fa - 4, ha - 0
                    fa #(.T(T)) fa72(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][5]}));
                    fa #(.T(T)) fa73(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][6]}));
                    fa #(.T(T)) fa74(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][7]}));
                    fa #(.T(T)) fa75(.i(s1[w][11:9]),.o({s2[w+1][3],s2[w][8]}));
                    assign s2[w][18:9] = s1[w][21:12];
                end
                42:
                begin
                    // fa - 3, ha - 0
                    fa #(.T(T)) fa76(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][4]}));
                    fa #(.T(T)) fa77(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][5]}));
                    fa #(.T(T)) fa78(.i(s1[w][8:6]),.o({s2[w+1][2],s2[w][6]}));
                    assign s2[w][18:7] = s1[w][20:9];
                end
                43:
                begin
                    // fa - 2, ha - 0
                    fa #(.T(T)) fa79(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][3]}));
                    fa #(.T(T)) fa80(.i(s1[w][5:3]),.o({s2[w+1][1],s2[w][4]}));
                    assign s2[w][18:5] = s1[w][19:6];
                end
                44:
                begin
                    // fa - 1, ha - 0
                    fa #(.T(T)) fa81(.i(s1[w][2:0]),.o({s2[w+1][0],s2[w][2]}));
                    assign s2[w][18:3] = s1[w][18:3];
                end
                45:
                begin
                    // carry
                    assign s2[w][18:1] = s1[w][17:0];
                end
                default:
                    assign s2[w] = s1[w];
            endcase 
        end
        // Stage 3 (Error could be here)
        // Max depth: 13 (12:0)
        for(w = 0;w <= 2*N-2;w = w+1)
        begin
            case(w)
                13:
                begin
                    // fa - 0, ha - 1
                    ha #(.T(T)) ha1(.i(s2[w][1:0]),.o({s3[w+1][0],s3[w][0]}));
                    assign s3[w][12:1] = s2[w][13:2];
                end
                14:
                begin
                    // fa - 1, ha - 1
                    fa #(.T(T)) fa1(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][1]}));
                    ha #(.T(T)) ha2(.i(s2[w][4:3]),.o({s3[w+1][1],s3[w][2]}));
                    assign s3[w][12:3] = s2[w][14:5];
                end
                15:
                begin
                    // fa - 2, ha - 1
                    fa #(.T(T)) fa2(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][2]}));
                    fa #(.T(T)) fa3(.i(s2[w][5:3]),.o({s3[w+1][1],s3[w][3]}));
                    ha #(.T(T)) ha3(.i(s2[w][7:6]),.o({s3[w+1][2],s3[w][4]}));
                    assign s3[w][12:5] = s2[w][15:8];
                end
                16:
                begin
                    // fa - 3, ha - 1
                    fa #(.T(T)) fa4(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][3]}));
                    fa #(.T(T)) fa5(.i(s2[w][5:3]),.o({s3[w+1][1],s3[w][4]}));
                    fa #(.T(T)) fa6(.i(s2[w][8:6]),.o({s3[w+1][2],s3[w][5]}));
                    ha #(.T(T)) ha4(.i(s2[w][10:9]),.o({s3[w+1][3],s3[w][6]}));
                    assign s3[w][12:7] = s2[w][16:11];
                end
                17:
                begin
                    // fa - 4, ha - 1
                    fa #(.T(T)) fa7(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][4]}));
                    fa #(.T(T)) fa8(.i(s2[w][5:3]),.o({s3[w+1][1],s3[w][5]}));
                    fa #(.T(T)) fa9(.i(s2[w][8:6]),.o({s3[w+1][2],s3[w][6]}));
                    fa #(.T(T)) fa10(.i(s2[w][11:9]),.o({s3[w+1][3],s3[w][7]}));
                    ha #(.T(T)) ha5(.i(s2[w][13:12]),.o({s3[w+1][4],s3[w][8]}));
                    assign s3[w][12:9] = s2[w][17:14];
                end
                18:
                begin
                    // fa - 5, ha - 1
                    fa #(.T(T)) fa11(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][5]}));
                    fa #(.T(T)) fa12(.i(s2[w][5:3]),.o({s3[w+1][1],s3[w][6]}));
                    fa #(.T(T)) fa13(.i(s2[w][8:6]),.o({s3[w+1][2],s3[w][7]}));
                    fa #(.T(T)) fa14(.i(s2[w][11:9]),.o({s3[w+1][3],s3[w][8]}));
                    fa #(.T(T)) fa15(.i(s2[w][14:12]),.o({s3[w+1][4],s3[w][9]}));
                    ha #(.T(T)) ha6(.i(s2[w][16:15]),.o({s3[w+1][5],s3[w][10]}));
                    assign s3[w][12:11] = s2[w][18:17];
                end
                19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45:
                begin
                    // fa - 6, ha - 0
                    fa #(.T(T)) fa16(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][6]}));
                    fa #(.T(T)) fa17(.i(s2[w][5:3]),.o({s3[w+1][1],s3[w][7]}));
                    fa #(.T(T)) fa18(.i(s2[w][8:6]),.o({s3[w+1][2],s3[w][8]}));
                    fa #(.T(T)) fa19(.i(s2[w][11:9]),.o({s3[w+1][3],s3[w][9]}));
                    fa #(.T(T)) fa20(.i(s2[w][14:12]),.o({s3[w+1][4],s3[w][10]}));
                    fa #(.T(T)) fa21(.i(s2[w][17:15]),.o({s3[w+1][5],s3[w][11]}));
                    assign s3[w][12] = s2[w][18];
                end
                46:
                begin
                    // fa - 5, ha - 0
                    fa #(.T(T)) fa22(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][6]}));
                    fa #(.T(T)) fa23(.i(s2[w][5:3]),.o({s3[w+1][1],s3[w][7]}));
                    fa #(.T(T)) fa24(.i(s2[w][8:6]),.o({s3[w+1][2],s3[w][8]}));
                    fa #(.T(T)) fa25(.i(s2[w][11:9]),.o({s3[w+1][3],s3[w][9]}));
                    fa #(.T(T)) fa26(.i(s2[w][14:12]),.o({s3[w+1][4],s3[w][10]}));
                    assign s3[w][12:11] = s2[w][16:15];
                end
                47:
                begin
                    // fa - 4, ha - 0
                    fa #(.T(T)) fa27(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][5]}));
                    fa #(.T(T)) fa28(.i(s2[w][5:3]),.o({s3[w+1][1],s3[w][6]}));
                    fa #(.T(T)) fa29(.i(s2[w][8:6]),.o({s3[w+1][2],s3[w][7]}));
                    fa #(.T(T)) fa30(.i(s2[w][11:9]),.o({s3[w+1][3],s3[w][8]}));
                    assign s3[w][12:9] = s2[w][15:12];
                end
                48:
                begin
                    // fa - 3, ha - 0
                    fa #(.T(T)) fa31(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][4]}));
                    fa #(.T(T)) fa32(.i(s2[w][5:3]),.o({s3[w+1][1],s3[w][5]}));
                    fa #(.T(T)) fa33(.i(s2[w][8:6]),.o({s3[w+1][2],s3[w][6]}));
                    assign s3[w][12:7] = s2[w][14:9];
                end
                49:
                begin
                    // fa - 2, ha - 0
                    fa #(.T(T)) fa34(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][3]}));
                    fa #(.T(T)) fa35(.i(s2[w][5:3]),.o({s3[w+1][1],s3[w][4]}));
                    assign s3[w][12:5] = s2[w][13:6];
                end
                50:
                begin
                    // fa - 1, ha - 0
                    fa #(.T(T)) fa36(.i(s2[w][2:0]),.o({s3[w+1][0],s3[w][2]}));
                    assign s3[w][12:3] = s2[w][12:3];
                end
                51:
                begin
                    // carry
                    assign s3[w][12:1] = s2[w][11:0];
                end
                default:
                    assign s3[w] = s2[w];
            endcase 
        end
        // Stage 4
        // Max depth: 9 (8:0)
        for(w = 0;w <= 2*N-2;w = w+1)
        begin
            case(w)
                9:
                begin
                    // fa - 0, ha - 1
                    ha #(.T(T)) ha1(.i(s3[w][1:0]),.o({s4[w+1][0],s4[w][0]}));
                    assign s4[w][8:1] = s3[w][9:2];
                end
                10:
                begin
                    // fa - 1, ha - 1
                    fa #(.T(T)) fa1(.i(s3[w][2:0]),.o({s4[w+1][0],s4[w][1]}));
                    ha #(.T(T)) ha2(.i(s3[w][4:3]),.o({s4[w+1][1],s4[w][2]}));
                    assign s4[w][8:3] = s3[w][10:5];
                end
                11:
                begin
                    // fa - 2, ha - 1
                    fa #(.T(T)) fa2(.i(s3[w][2:0]),.o({s4[w+1][0],s4[w][2]}));
                    fa #(.T(T)) fa3(.i(s3[w][5:3]),.o({s4[w+1][1],s4[w][3]}));
                    ha #(.T(T)) ha3(.i(s3[w][7:6]),.o({s4[w+1][2],s4[w][4]}));
                    assign s4[w][8:5] = s3[w][11:8];
                end
                12:
                begin
                    // fa - 3, ha - 1
                    fa #(.T(T)) fa4(.i(s3[w][2:0]),.o({s4[w+1][0],s4[w][3]}));
                    fa #(.T(T)) fa5(.i(s3[w][5:3]),.o({s4[w+1][1],s4[w][4]}));
                    fa #(.T(T)) fa6(.i(s3[w][8:6]),.o({s4[w+1][2],s4[w][5]}));
                    ha #(.T(T)) ha4(.i(s3[w][10:9]),.o({s4[w+1][3],s4[w][6]}));
                    assign s4[w][8:7] = s3[w][12:11];
                end
                13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51:
                begin
                    // fa - 4, ha - 0
                    fa #(.T(T)) fa7(.i(s3[w][2:0]),.o({s4[w+1][0],s4[w][4]}));
                    fa #(.T(T)) fa8(.i(s3[w][5:3]),.o({s4[w+1][1],s4[w][5]}));
                    fa #(.T(T)) fa9(.i(s3[w][8:6]),.o({s4[w+1][2],s4[w][6]}));
                    fa #(.T(T)) fa10(.i(s3[w][11:9]),.o({s4[w+1][3],s4[w][7]}));
                    assign s4[w][8] = s3[w][12];
                end
                52:
                begin
                    // fa - 3, ha - 0
                    fa #(.T(T)) fa11(.i(s3[w][2:0]),.o({s4[w+1][0],s4[w][4]}));
                    fa #(.T(T)) fa12(.i(s3[w][5:3]),.o({s4[w+1][1],s4[w][5]}));
                    fa #(.T(T)) fa13(.i(s3[w][8:6]),.o({s4[w+1][2],s4[w][6]}));
                    assign s4[w][8:7] = s3[w][10:9];
                end
                53:
                begin
                    // fa - 2, ha - 0
                    fa #(.T(T)) fa14(.i(s3[w][2:0]),.o({s4[w+1][0],s4[w][3]}));
                    fa #(.T(T)) fa15(.i(s3[w][5:3]),.o({s4[w+1][1],s4[w][4]}));
                    assign s4[w][8:5] = s3[w][9:6];
                end
                54:
                begin
                    // fa - 1, ha - 0
                    fa #(.T(T)) fa16(.i(s3[w][2:0]),.o({s4[w+1][0],s4[w][2]}));
                    assign s4[w][8:3] = s3[w][8:3];
                end
                55:
                begin
                    // carry
                    assign s4[w][8:1] = s3[w][7:0];
                end
                default:
                    assign s4[w] = s3[w];
            endcase 
        end
        // Stage 5
        // Max depth: 6 (5:0)
        for(w = 0;w <= 2*N-2;w = w+1)
        begin
            case(w)
                6:
                begin 
                    // fa - 0, ha - 1
                    ha #(.T(T)) ha1(.i(s4[w][1:0]),.o({s5[w+1][0],s5[w][0]}));
                    assign s5[w][5:1] = s4[w][6:2];
                end
                7:
                begin
                    // fa - 1, ha - 1
                    fa #(.T(T)) fa1(.i(s4[w][2:0]),.o({s5[w+1][0],s5[w][1]}));
                    ha #(.T(T)) ha2(.i(s4[w][4:3]),.o({s5[w+1][1],s5[w][2]}));
                    assign s5[w][5:3] = s4[w][7:5];
                end
                8:
                begin
                    // fa - 2, ha - 1
                    fa #(.T(T)) fa2(.i(s4[w][2:0]),.o({s5[w+1][0],s5[w][2]}));
                    fa #(.T(T)) fa3(.i(s4[w][5:3]),.o({s5[w+1][1],s5[w][3]}));
                    ha #(.T(T)) ha3(.i(s4[w][7:6]),.o({s5[w+1][2],s5[w][4]}));
                    assign s5[w][5] = s4[w][8];
                end
                9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55:
                begin
                    // fa - 3, ha - 0
                    fa #(.T(T)) fa4(.i(s4[w][2:0]),.o({s5[w+1][0],s5[w][3]}));
                    fa #(.T(T)) fa5(.i(s4[w][5:3]),.o({s5[w+1][1],s5[w][4]}));
                    fa #(.T(T)) fa6(.i(s4[w][8:6]),.o({s5[w+1][2],s5[w][5]}));
                end
                56:
                begin
                    // fa - 2, ha - 0
                    fa #(.T(T)) fa7(.i(s4[w][2:0]),.o({s5[w+1][0],s5[w][3]}));
                    fa #(.T(T)) fa8(.i(s4[w][5:3]),.o({s5[w+1][1],s5[w][4]}));
                    assign s5[w][5] = s4[w][6];
                end
                57:
                begin
                    // fa - 1, ha - 0
                    fa #(.T(T)) fa9(.i(s4[w][2:0]),.o({s5[w+1][0],s5[w][2]}));
                    assign s5[w][5:3] = s4[w][5:3];
                end
                58:
                begin
                    // carry
                    assign s5[w][5:1] = s4[w][4:0];
                end
                default:
                    assign s5[w] = s4[w];
            endcase 
        end
        // Stage 6
        // Max depth: 4 (3:0)
        for(w = 0;w <= 2*N-2;w = w+1)
        begin
            case(w)
                4:
                begin 
                    // fa - 0, ha - 1
                    ha #(.T(T)) ha1(.i(s5[w][1:0]),.o({s6[w+1][0],s6[w][0]}));
                    assign s6[w][3:1] = s5[w][4:2];
                end
                5:
                begin
                    // fa - 1, ha - 1
                    fa #(.T(T)) fa1(.i(s5[w][2:0]),.o({s6[w+1][0],s6[w][1]}));
                    ha #(.T(T)) ha2(.i(s5[w][4:3]),.o({s6[w+1][1],s6[w][2]}));
                    assign s6[w][3] = s5[w][5];
                end
                6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58:
                begin
                    // fa - 2, ha - 0
                    fa #(.T(T)) fa4(.i(s5[w][2:0]),.o({s6[w+1][0],s6[w][2]}));
                    fa #(.T(T)) fa5(.i(s5[w][5:3]),.o({s6[w+1][1],s6[w][3]}));
                end
                59:
                begin
                    // fa - 1, ha - 0
                    fa #(.T(T)) fa6(.i(s5[w][2:0]),.o({s6[w+1][0],s6[w][2]}));
                    assign s6[w][3] = s5[w][3];
                end
                60:
                begin
                    // carry
                    assign s6[w][3:1] = s5[w][2:0];
                end
                default:
                    assign s6[w] = s5[w];
            endcase 
        end
        // Stage 7
        // Max depth: 3 (2:0)
        for(w = 0;w <= 2*N-2;w = w+1)
        begin
            case(w)
                3:
                begin 
                    // fa - 0, ha - 1
                    ha #(.T(T)) ha1(.i(s6[w][1:0]),.o({s7[w+1][0],s7[w][0]}));
                    assign s7[w][2:1] = s6[w][3:2];
                end
                4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60:
                begin
                    // fa - 1, ha - 0
                    fa #(.T(T)) fa1(.i(s6[w][2:0]),.o({s7[w+1][0],s7[w][1]}));
                    assign s7[w][2] = s6[w][3];
                end
                61:
                begin
                    // fa - carry
                    assign s7[w][2:1] = s6[w][1:0];
                end
                default:
                    assign s7[w] = s6[w];
            endcase 
        end
        // Stage 8
        // Max depth: 2 (1:0)
        for(w = 0;w <= 2*N-2;w = w+1)
        begin
            case(w)
                2:
                begin 
                    // fa - 0, ha - 1
                    ha #(.T(T)) ha1(.i(s7[w][1:0]),.o({s8[w+1][0],s8[w][0]}));
                    assign s8[w][1] = s7[w][2];
                end
                3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61:
                begin
                    // fa - 1, ha - 0
                    fa #(.T(T)) fa1(.i(s7[w][2:0]),.o({s8[w+1][0],s8[w][1]}));
                end
                62:
                begin
                    // fa - carry
                    assign s8[w][1] = s7[w][0];
                end
                default:
                    assign s8[w] = s7[w];
            endcase 
        end
    endgenerate
    add32 #(.T(T)) add0(
        .a({s8[31][0],s8[30][0],s8[29][0],s8[28][0],s8[27][0],s8[26][0],s8[25][0],s8[24][0],s8[23][0],s8[22][0],s8[21][0],s8[20][0],s8[19][0],s8[18][0],s8[17][0],s8[16][0],s8[15][0],s8[14][0],s8[13][0],s8[12][0],s8[11][0],s8[10][0],s8[9][0],s8[8][0],s8[7][0],s8[6][0],s8[5][0],s8[4][0],s8[3][0],s8[2][0],s8[1][0],s8[0][0]}),
        .b({s8[31][1],s8[30][1],s8[29][1],s8[28][1],s8[27][1],s8[26][1],s8[25][1],s8[24][1],s8[23][1],s8[22][1],s8[21][1],s8[20][1],s8[19][1],s8[18][1],s8[17][1],s8[16][1],s8[15][1],s8[14][1],s8[13][1],s8[12][1],s8[11][1],s8[10][1],s8[9][1],s8[8][1],s8[7][1],s8[6][1],s8[5][1],s8[4][1],s8[3][1],s8[2][1],s8[1][1],1'b0}),
        .c_1(1'b0),
        .s(lo_),
        .c31(c)
    );
    add32 #(.T(T)) add1(
        .a({1'b0, s8[62][0],s8[61][0],s8[60][0],s8[59][0],s8[58][0],s8[57][0],s8[56][0],s8[55][0],s8[54][0],s8[53][0],s8[52][0],s8[51][0],s8[50][0],s8[49][0],s8[48][0],s8[47][0],s8[46][0],s8[45][0],s8[44][0],s8[43][0],s8[42][0],s8[41][0],s8[40][0],s8[39][0],s8[38][0],s8[37][0],s8[36][0],s8[35][0],s8[34][0],s8[33][0],s8[32][0]}),
        .b({1'b0, s8[62][1],s8[61][1],s8[60][1],s8[59][1],s8[58][1],s8[57][1],s8[56][1],s8[55][1],s8[54][1],s8[53][1],s8[52][1],s8[51][1],s8[50][1],s8[49][1],s8[48][1],s8[47][1],s8[46][1],s8[45][1],s8[44][1],s8[43][1],s8[42][1],s8[41][1],s8[40][1],s8[39][1],s8[38][1],s8[37][1],s8[36][1],s8[35][1],s8[34][1],s8[33][1],s8[32][1]}),
        .c_1(c),
        .s(hi_)
    );
    add32 #(.T(T)) add2(
        .a(lo__),
        .b(32'h00000000),
        .c_1(prod_comp),
        .s(lo),
        .c31(c_)
    );
    add32 #(.T(T)) add3(
        .a(hi__),
        .b(32'h00000000),
        .c_1(c_),
        .s(hi)
    );
endmodule