module datapath #(parameter T = 32) (
    input clk
);