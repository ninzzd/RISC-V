module alu(
    input [31:0] a,
    input [31:0] b,
    input alu_ctrl,
    output [31:0] lo,
    output [31:0] hi
);
endmodule