module l1_data_cache(
    input [31:0] addr,
    input WE,
    input [31:0] wd,
    output [31:0] rd;
);
endmodule 