module l1_instr_cache #(parameter size = 8192, parameter Clen = $clog2(size))(
    
);
endmodule