module qru(
    input [31:0] a,
    input [31:0] b,
    input [1:0] divctl,
    output [31:0] res
);

endmodule