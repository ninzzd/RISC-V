module l1_data_cache(

);
endmodule 