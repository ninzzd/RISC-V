module shift_right32(
    input [31:0] inp,
    input [4:0] shamt,
    input mode, // mode: 0 => srl, 1 -> sra
    output [31:0] res
);
    wire s;
    wire [31:0] in0;
    wire [31:0] in1;
    wire [31:0] in2;
    wire [31:0] in3;
    wire [31:0] in4;
    wire [31:0] in5;
    wire [31:0] in6;
    wire [31:0] in7;
    wire [31:0] in8;
    wire [31:0] in9;
    wire [31:0] in10;
    wire [31:0] in11;
    wire [31:0] in12;
    wire [31:0] in13;
    wire [31:0] in14;
    wire [31:0] in15;
    wire [31:0] in16;
    wire [31:0] in17;
    wire [31:0] in18;
    wire [31:0] in19;
    wire [31:0] in20;
    wire [31:0] in21;
    wire [31:0] in22;
    wire [31:0] in23;
    wire [31:0] in24;
    wire [31:0] in25;
    wire [31:0] in26;
    wire [31:0] in27;
    wire [31:0] in28;
    wire [31:0] in29;
    wire [31:0] in30;
    wire [31:0] in31;

    assign s = mode&inp[31];
    assign in0  = inp;
    assign in1  = {s,inp[31:1]};
    assign in2  = {{2{s}},inp[31:2]};
    assign in3  = {{3{s}},inp[31:3]};
    assign in4  = {{4{s}},inp[31:4]};
    assign in5  = {{5{s}},inp[31:5]};
    assign in6  = {{6{s}},inp[31:6]};
    assign in7  = {{7{s}},inp[31:7]};
    assign in8  = {{8{s}},inp[31:8]};
    assign in9  = {{9{s}},inp[31:9]};
    assign in10 = {{10{s}},inp[31:10]};
    assign in11 = {{11{s}},inp[31:11]};
    assign in12 = {{12{s}},inp[31:12]};
    assign in13 = {{13{s}},inp[31:13]};
    assign in14 = {{14{s}},inp[31:14]};
    assign in15 = {{15{s}},inp[31:15]};
    assign in16 = {{16{s}},inp[31:16]};
    assign in17 = {{17{s}},inp[31:17]};
    assign in18 = {{18{s}},inp[31:18]};
    assign in19 = {{19{s}},inp[31:19]};
    assign in20 = {{20{s}},inp[31:20]};
    assign in21 = {{21{s}},inp[31:21]};
    assign in22 = {{22{s}},inp[31:22]};
    assign in23 = {{23{s}},inp[31:23]};
    assign in24 = {{24{s}},inp[31:24]};
    assign in25 = {{25{s}},inp[31:25]};
    assign in26 = {{26{s}},inp[31:26]};
    assign in27 = {{27{s}},inp[31:27]};
    assign in28 = {{28{s}},inp[31:28]};
    assign in29 = {{29{s}},inp[31:29]};
    assign in30 = {{30{s}},inp[31:30]};
    assign in31 = {{30{s}},inp[31]};
    
    mux32t1 m0(.in(in0),.sel(shamt),.out(res[0]));
    mux32t1 m1(.in(in1),.sel(shamt),.out(res[1]));
    mux32t1 m2(.in(in2),.sel(shamt),.out(res[2]));
    mux32t1 m3(.in(in3),.sel(shamt),.out(res[3]));
    mux32t1 m4(.in(in4),.sel(shamt),.out(res[4]));
    mux32t1 m5(.in(in5),.sel(shamt),.out(res[5]));
    mux32t1 m6(.in(in6),.sel(shamt),.out(res[6]));
    mux32t1 m7(.in(in7),.sel(shamt),.out(res[7]));
    mux32t1 m8(.in(in8),.sel(shamt),.out(res[8]));
    mux32t1 m9(.in(in9),.sel(shamt),.out(res[9]));
    mux32t1 m10(.in(in10),.sel(shamt),.out(res[10]));
    mux32t1 m11(.in(in11),.sel(shamt),.out(res[11]));
    mux32t1 m12(.in(in12),.sel(shamt),.out(res[12]));
    mux32t1 m13(.in(in13),.sel(shamt),.out(res[13]));
    mux32t1 m14(.in(in14),.sel(shamt),.out(res[14]));
    mux32t1 m15(.in(in15),.sel(shamt),.out(res[15]));
    mux32t1 m16(.in(in16),.sel(shamt),.out(res[16]));
    mux32t1 m17(.in(in17),.sel(shamt),.out(res[17]));
    mux32t1 m18(.in(in18),.sel(shamt),.out(res[18]));
    mux32t1 m19(.in(in19),.sel(shamt),.out(res[19]));
    mux32t1 m20(.in(in20),.sel(shamt),.out(res[20]));
    mux32t1 m21(.in(in21),.sel(shamt),.out(res[21]));
    mux32t1 m22(.in(in22),.sel(shamt),.out(res[22]));
    mux32t1 m23(.in(in23),.sel(shamt),.out(res[23]));
    mux32t1 m24(.in(in24),.sel(shamt),.out(res[24]));
    mux32t1 m25(.in(in25),.sel(shamt),.out(res[25]));
    mux32t1 m26(.in(in26),.sel(shamt),.out(res[26]));
    mux32t1 m27(.in(in27),.sel(shamt),.out(res[27]));
    mux32t1 m28(.in(in28),.sel(shamt),.out(res[28]));
    mux32t1 m29(.in(in29),.sel(shamt),.out(res[29]));
    mux32t1 m30(.in(in30),.sel(shamt),.out(res[30]));
    mux32t1 m31(.in(in31),.sel(shamt),.out(res[31]));
endmodule