module shift32(
    input [31:0] operand,
    input [4:0] shamt,
    input mode,
    output [31:0] res
);

endmodule