`timescale 1ns/1ps
module riscv_tb;
    // Testbench code for RISC-V processor would go here
endmodule
