module risc_v #(parameter T = 0.000)(

);
endmodule
