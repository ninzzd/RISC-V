module shift_left32(
    input [31:0] inp,
    input [4:0] shamt,
    input mode,
    output [31:0] res
);
    wire [31:0] in0;
    wire [31:0] in1;
    wire [31:0] in2;
    wire [31:0] in3;
    wire [31:0] in4;
    wire [31:0] in5;
    wire [31:0] in6;
    wire [31:0] in7;
    wire [31:0] in8;
    wire [31:0] in9;
    wire [31:0] in10;
    wire [31:0] in11;
    wire [31:0] in12;
    wire [31:0] in13;
    wire [31:0] in14;
    wire [31:0] in15;
    wire [31:0] in16;
    wire [31:0] in17;
    wire [31:0] in18;
    wire [31:0] in19;
    wire [31:0] in20;
    wire [31:0] in21;
    wire [31:0] in22;
    wire [31:0] in23;
    wire [31:0] in24;
    wire [31:0] in25;
    wire [31:0] in26;
    wire [31:0] in27;
    wire [31:0] in28;
    wire [31:0] in29;
    wire [31:0] in30;
    wire [31:0] in31;

    assign in0  = {{31{1'b0}},{inp[0]}};
    assign in1  = {{30{1'b0}},{inp[0],inp[1]}};
    assign in2  = {{29{1'b0}},{inp[0],inp[1],inp[2]}};
    assign in3  = {{28{1'b0}},{inp[0],inp[1],inp[2],inp[3]}};
    assign in4  = {{27{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4]}};
    assign in5  = {{26{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5]}};
    assign in6  = {{25{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6]}};
    assign in7  = {{24{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7]}};
    assign in8  = {{23{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8]}};
    assign in9  = {{22{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9]}};
    assign in10 = {{21{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10]}};
    assign in11 = {{20{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11]}};
    assign in12 = {{19{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12]}};
    assign in13 = {{18{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13]}};
    assign in14 = {{17{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14]}};
    assign in15 = {{16{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15]}};
    assign in16 = {{15{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16]}};
    assign in17 = {{14{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17]}};
    assign in18 = {{13{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18]}};
    assign in19 = {{12{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19]}};
    assign in20 = {{11{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20]}};
    assign in21 = {{10{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21]}};
    assign in22 = {{9{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21],inp[22]}};
    assign in23 = {{8{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21],inp[22],inp[23]}};
    assign in24 = {{7{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21],inp[22],inp[23],inp[24]}};
    assign in25 = {{6{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21],inp[22],inp[23],inp[24],inp[25]}};
    assign in26 = {{5{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21],inp[22],inp[23],inp[24],inp[25],inp[26]}};
    assign in27 = {{4{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21],inp[22],inp[23],inp[24],inp[25],inp[26],inp[27]}};
    assign in28 = {{3{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21],inp[22],inp[23],inp[24],inp[25],inp[26],inp[27],inp[28]}};
    assign in29 = {{2{1'b0}},{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21],inp[22],inp[23],inp[24],inp[25],inp[26],inp[27],inp[28],inp[29]}};
    assign in30 = {1'b0,{inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21],inp[22],inp[23],inp[24],inp[25],inp[26],inp[27],inp[28],inp[29],inp[30]}};
    assign in31 = {inp[0],inp[1],inp[2],inp[3],inp[4],inp[5],inp[6],inp[7],inp[8],inp[9],inp[10],inp[11],inp[12],inp[13],inp[14],inp[15],inp[16],inp[17],inp[18],inp[19],inp[20],inp[21],inp[22],inp[23],inp[24],inp[25],inp[26],inp[27],inp[28],inp[29],inp[30],inp[31]};
    
    mux32t1 m0(.in(in0),.sel(shamt),.out(res[0]));
    mux32t1 m1(.in(in1),.sel(shamt),.out(res[1]));
    mux32t1 m2(.in(in2),.sel(shamt),.out(res[2]));
    mux32t1 m3(.in(in3),.sel(shamt),.out(res[3]));
    mux32t1 m4(.in(in4),.sel(shamt),.out(res[4]));
    mux32t1 m5(.in(in5),.sel(shamt),.out(res[5]));
    mux32t1 m6(.in(in6),.sel(shamt),.out(res[6]));
    mux32t1 m7(.in(in7),.sel(shamt),.out(res[7]));
    mux32t1 m8(.in(in8),.sel(shamt),.out(res[8]));
    mux32t1 m9(.in(in9),.sel(shamt),.out(res[9]));
    mux32t1 m10(.in(in10),.sel(shamt),.out(res[10]));
    mux32t1 m11(.in(in11),.sel(shamt),.out(res[11]));
    mux32t1 m12(.in(in12),.sel(shamt),.out(res[12]));
    mux32t1 m13(.in(in13),.sel(shamt),.out(res[13]));
    mux32t1 m14(.in(in14),.sel(shamt),.out(res[14]));
    mux32t1 m15(.in(in15),.sel(shamt),.out(res[15]));
    mux32t1 m16(.in(in16),.sel(shamt),.out(res[16]));
    mux32t1 m17(.in(in17),.sel(shamt),.out(res[17]));
    mux32t1 m18(.in(in18),.sel(shamt),.out(res[18]));
    mux32t1 m19(.in(in19),.sel(shamt),.out(res[19]));
    mux32t1 m20(.in(in20),.sel(shamt),.out(res[20]));
    mux32t1 m21(.in(in21),.sel(shamt),.out(res[21]));
    mux32t1 m22(.in(in22),.sel(shamt),.out(res[22]));
    mux32t1 m23(.in(in23),.sel(shamt),.out(res[23]));
    mux32t1 m24(.in(in24),.sel(shamt),.out(res[24]));
    mux32t1 m25(.in(in25),.sel(shamt),.out(res[25]));
    mux32t1 m26(.in(in26),.sel(shamt),.out(res[26]));
    mux32t1 m27(.in(in27),.sel(shamt),.out(res[27]));
    mux32t1 m28(.in(in28),.sel(shamt),.out(res[28]));
    mux32t1 m29(.in(in29),.sel(shamt),.out(res[29]));
    mux32t1 m30(.in(in30),.sel(shamt),.out(res[30]));
    mux32t1 m31(.in(in31),.sel(shamt),.out(res[31]));
endmodule